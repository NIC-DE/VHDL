--libr