-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
-- CREATED		"Wed Sep 16 20:01:52 2020"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY decoder IS 
	PORT
	(
		CLK :  IN  STD_LOGIC;
		CE :  IN  STD_LOGIC;
		CLR :  IN  STD_LOGIC;
		Carry :  IN  STD_LOGIC;
		Zero :  IN  STD_LOGIC;
		IR :  IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		EN_PC :  OUT  STD_LOGIC;
		EN_DA :  OUT  STD_LOGIC;
		EN_IN :  OUT  STD_LOGIC;
		MUXC :  OUT  STD_LOGIC;
		MUXB :  OUT  STD_LOGIC;
		MUXA :  OUT  STD_LOGIC;
		ALU_S4 :  OUT  STD_LOGIC;
		ALU_S3 :  OUT  STD_LOGIC;
		ALU_S2 :  OUT  STD_LOGIC;
		ALU_S0 :  OUT  STD_LOGIC;
		RAM :  OUT  STD_LOGIC;
		ALU_S1 :  OUT  STD_LOGIC
	);
END decoder;

ARCHITECTURE bdf_type OF decoder IS 

COMPONENT sequence_generator
	PORT(CLK : IN STD_LOGIC;
		 CE : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 FETCH : OUT STD_LOGIC;
		 DECODE : OUT STD_LOGIC;
		 EXECUTE : OUT STD_LOGIC;
		 INCREMENT : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT status_register
	PORT(Carry : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 Zero : IN STD_LOGIC;
		 ADD : IN STD_LOGIC;
		 SUB : IN STD_LOGIC;
		 BITAND : IN STD_LOGIC;
		 CARRY_REG : OUT STD_LOGIC;
		 ZERO_REG : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT instruction_decoder_full
	PORT(DECODE : IN STD_LOGIC;
		 EXECUTE : IN STD_LOGIC;
		 IR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		 INPUT : OUT STD_LOGIC;
		 OUTPUT : OUT STD_LOGIC;
		 LOAD : OUT STD_LOGIC;
		 ADD : OUT STD_LOGIC;
		 JUMPZ : OUT STD_LOGIC;
		 JUMP : OUT STD_LOGIC;
		 JUMPNZ : OUT STD_LOGIC;
		 JUMPC : OUT STD_LOGIC;
		 JUMPNC : OUT STD_LOGIC;
		 SUB : OUT STD_LOGIC;
		 BITAND : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT jump_detector
	PORT(INCREMENT : IN STD_LOGIC;
		 EXECUTE : IN STD_LOGIC;
		 ZERO_REG : IN STD_LOGIC;
		 CARRY_REG : IN STD_LOGIC;
		 JUMPZ : IN STD_LOGIC;
		 JUMPNZ : IN STD_LOGIC;
		 JUMPC : IN STD_LOGIC;
		 JUMPNC : IN STD_LOGIC;
		 JUMP : IN STD_LOGIC;
		 CLK : IN STD_LOGIC;
		 CLR : IN STD_LOGIC;
		 EN_PC : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_65 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_66 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_67 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_68 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_69 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_70 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_52 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_53 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_54 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_12 <= '0';
SYNTHESIZED_WIRE_29 <= '0';



b2v_inst : sequence_generator
PORT MAP(CLK => CLK,
		 CE => CE,
		 CLR => CLR,
		 FETCH => SYNTHESIZED_WIRE_52,
		 DECODE => SYNTHESIZED_WIRE_41,
		 EXECUTE => SYNTHESIZED_WIRE_58,
		 INCREMENT => SYNTHESIZED_WIRE_64);

ALU_S3 <= SYNTHESIZED_WIRE_57;


ALU_S2 <= SYNTHESIZED_WIRE_1;


ALU_S1 <= SYNTHESIZED_WIRE_2;


ALU_S0 <= SYNTHESIZED_WIRE_3;


RAM <= SYNTHESIZED_WIRE_4;



SYNTHESIZED_WIRE_40 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_6;


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_60 OR SYNTHESIZED_WIRE_61 OR SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_12;



SYNTHESIZED_WIRE_53 <= SYNTHESIZED_WIRE_63 OR SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_54 <= SYNTHESIZED_WIRE_61 OR SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_60;


b2v_inst2 : status_register
PORT MAP(Carry => Carry,
		 CLK => CLK,
		 CLR => CLR,
		 Zero => Zero,
		 ADD => SYNTHESIZED_WIRE_60,
		 SUB => SYNTHESIZED_WIRE_57,
		 BITAND => SYNTHESIZED_WIRE_62,
		 CARRY_REG => SYNTHESIZED_WIRE_46,
		 ZERO_REG => SYNTHESIZED_WIRE_45);


SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_57 OR SYNTHESIZED_WIRE_64;


SYNTHESIZED_WIRE_70 <= SYNTHESIZED_WIRE_65 OR SYNTHESIZED_WIRE_66 OR SYNTHESIZED_WIRE_67 OR SYNTHESIZED_WIRE_68 OR SYNTHESIZED_WIRE_69 OR SYNTHESIZED_WIRE_29;



SYNTHESIZED_WIRE_2 <= SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_63 OR SYNTHESIZED_WIRE_61 OR SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_3 <= SYNTHESIZED_WIRE_70 OR SYNTHESIZED_WIRE_61 OR SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_4 <= SYNTHESIZED_WIRE_58 AND SYNTHESIZED_WIRE_63;

EN_DA <= SYNTHESIZED_WIRE_40;



b2v_inst3 : instruction_decoder_full
PORT MAP(DECODE => SYNTHESIZED_WIRE_41,
		 EXECUTE => SYNTHESIZED_WIRE_58,
		 IR => IR,
		 INPUT => SYNTHESIZED_WIRE_59,
		 OUTPUT => SYNTHESIZED_WIRE_63,
		 LOAD => SYNTHESIZED_WIRE_61,
		 ADD => SYNTHESIZED_WIRE_60,
		 JUMPZ => SYNTHESIZED_WIRE_65,
		 JUMP => SYNTHESIZED_WIRE_69,
		 JUMPNZ => SYNTHESIZED_WIRE_67,
		 JUMPC => SYNTHESIZED_WIRE_66,
		 JUMPNC => SYNTHESIZED_WIRE_68,
		 SUB => SYNTHESIZED_WIRE_57,
		 BITAND => SYNTHESIZED_WIRE_62);


b2v_inst4 : jump_detector
PORT MAP(INCREMENT => SYNTHESIZED_WIRE_64,
		 EXECUTE => SYNTHESIZED_WIRE_58,
		 ZERO_REG => SYNTHESIZED_WIRE_45,
		 CARRY_REG => SYNTHESIZED_WIRE_46,
		 JUMPZ => SYNTHESIZED_WIRE_65,
		 JUMPNZ => SYNTHESIZED_WIRE_67,
		 JUMPC => SYNTHESIZED_WIRE_66,
		 JUMPNC => SYNTHESIZED_WIRE_68,
		 JUMP => SYNTHESIZED_WIRE_69,
		 CLK => CLK,
		 CLR => CLR,
		 EN_PC => EN_PC);

EN_IN <= SYNTHESIZED_WIRE_52;


MUXC <= SYNTHESIZED_WIRE_53;


MUXB <= SYNTHESIZED_WIRE_54;


MUXA <= SYNTHESIZED_WIRE_64;


ALU_S4 <= SYNTHESIZED_WIRE_64;



END bdf_type;